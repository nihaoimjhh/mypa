//Generate the verilog at 2024-08-18T18:18:20
module top (
BTN,
LD,
SW1,
SW2
);

input [2:0] BTN ;
output [6:0] LD ;
input [3:0] SW1 ;
input [3:0] SW2 ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire \add3/_00_ ;
wire \add3/_01_ ;
wire \add3/_02_ ;
wire \add3/_03_ ;
wire \add3/_04_ ;
wire \add3/_05_ ;
wire \add3/_06_ ;
wire \add3/_07_ ;
wire \add3/cout1 ;
wire \add3/cout2 ;
wire \add3/cout3 ;
wire \add3/cout4 ;
wire \add3/s0 ;
wire \add3/s1 ;
wire \add3/s2 ;
wire \add3/s3 ;
wire \add3/insert_0/_00_ ;
wire \add3/insert_0/_01_ ;
wire \add3/insert_0/_02_ ;
wire \add3/insert_0/_03_ ;
wire \add3/insert_0/_04_ ;
wire \add3/insert_0/_05_ ;
wire \add3/insert_0/_06_ ;
wire \add3/insert_0/_07_ ;
wire \add3/insert_1/_00_ ;
wire \add3/insert_1/_01_ ;
wire \add3/insert_1/_02_ ;
wire \add3/insert_1/_03_ ;
wire \add3/insert_1/_04_ ;
wire \add3/insert_1/_05_ ;
wire \add3/insert_1/_06_ ;
wire \add3/insert_1/_07_ ;
wire \add3/insert_2/_00_ ;
wire \add3/insert_2/_01_ ;
wire \add3/insert_2/_02_ ;
wire \add3/insert_2/_03_ ;
wire \add3/insert_2/_04_ ;
wire \add3/insert_2/_05_ ;
wire \add3/insert_2/_06_ ;
wire \add3/insert_2/_07_ ;
wire \add3/insert_3/_00_ ;
wire \add3/insert_3/_01_ ;
wire \add3/insert_3/_02_ ;
wire \add3/insert_3/_03_ ;
wire \add3/insert_3/_04_ ;
wire \add3/insert_3/_05_ ;
wire \add3/insert_3/_06_ ;
wire \add3/insert_3/_07_ ;
wire \and3/_00_ ;
wire \and3/_01_ ;
wire \and3/_02_ ;
wire \and3/_03_ ;
wire \and3/_04_ ;
wire \and3/_05_ ;
wire \and3/_06_ ;
wire \and3/_07_ ;
wire \and3/_08_ ;
wire \and3/_09_ ;
wire \and3/_10_ ;
wire \and3/_11_ ;
wire \and3/_12_ ;
wire \c3/_00_ ;
wire \c3/_01_ ;
wire \c3/_02_ ;
wire \c3/_03_ ;
wire \c3/_04_ ;
wire \c3/_05_ ;
wire \c3/_06_ ;
wire \c3/_07_ ;
wire \c3/_08_ ;
wire \c3/_09_ ;
wire \c3/_10_ ;
wire \c3/_11_ ;
wire \c3/_12_ ;
wire \c3/_13_ ;
wire \c3/_14_ ;
wire \c3/_15_ ;
wire \c3/_16_ ;
wire \c3/_17_ ;
wire \c3/_18_ ;
wire \c3/_19_ ;
wire \c3/_20_ ;
wire \c3/_21_ ;
wire \c3/eq0 ;
wire \eq3/_00_ ;
wire \eq3/_01_ ;
wire \eq3/_02_ ;
wire \eq3/_03_ ;
wire \eq3/_04_ ;
wire \eq3/_05_ ;
wire \eq3/_06_ ;
wire \eq3/_07_ ;
wire \eq3/_08_ ;
wire \eq3/_09_ ;
wire \eq3/eq0 ;
wire \not3/_00_ ;
wire \not3/_01_ ;
wire \not3/_02_ ;
wire \not3/_03_ ;
wire \not3/_04_ ;
wire \not3/_05_ ;
wire \not3/_06_ ;
wire \not3/_07_ ;
wire \not3/_08_ ;
wire \or3/_00_ ;
wire \or3/_01_ ;
wire \or3/_02_ ;
wire \or3/_03_ ;
wire \or3/_04_ ;
wire \or3/_05_ ;
wire \or3/_06_ ;
wire \or3/_07_ ;
wire \or3/_08_ ;
wire \or3/_09_ ;
wire \or3/_10_ ;
wire \or3/_11_ ;
wire \or3/_12_ ;
wire \sub3/_00_ ;
wire \sub3/_01_ ;
wire \sub3/_02_ ;
wire \sub3/_03_ ;
wire \sub3/_04_ ;
wire \sub3/_05_ ;
wire \sub3/_06_ ;
wire \sub3/insert_0/_00_ ;
wire \sub3/insert_0/_01_ ;
wire \sub3/insert_0/_02_ ;
wire \sub3/insert_0/_03_ ;
wire \sub3/insert_0/_04_ ;
wire \sub3/insert_0/_05_ ;
wire \sub3/insert_0/_06_ ;
wire \sub3/insert_0/_07_ ;
wire \sub3/insert_0/cout1 ;
wire \sub3/insert_0/cout2 ;
wire \sub3/insert_0/cout3 ;
wire \sub3/insert_0/cout4 ;
wire \sub3/insert_0/s0 ;
wire \sub3/insert_0/s1 ;
wire \sub3/insert_0/s2 ;
wire \sub3/insert_0/s3 ;
wire \sub3/insert_0/insert_0/_00_ ;
wire \sub3/insert_0/insert_0/_01_ ;
wire \sub3/insert_0/insert_0/_02_ ;
wire \sub3/insert_0/insert_0/_03_ ;
wire \sub3/insert_0/insert_0/_04_ ;
wire \sub3/insert_0/insert_0/_05_ ;
wire \sub3/insert_0/insert_0/_06_ ;
wire \sub3/insert_0/insert_0/_07_ ;
wire \sub3/insert_0/insert_1/_00_ ;
wire \sub3/insert_0/insert_1/_01_ ;
wire \sub3/insert_0/insert_1/_02_ ;
wire \sub3/insert_0/insert_1/_03_ ;
wire \sub3/insert_0/insert_1/_04_ ;
wire \sub3/insert_0/insert_1/_05_ ;
wire \sub3/insert_0/insert_1/_06_ ;
wire \sub3/insert_0/insert_1/_07_ ;
wire \sub3/insert_0/insert_2/_00_ ;
wire \sub3/insert_0/insert_2/_01_ ;
wire \sub3/insert_0/insert_2/_02_ ;
wire \sub3/insert_0/insert_2/_03_ ;
wire \sub3/insert_0/insert_2/_04_ ;
wire \sub3/insert_0/insert_2/_05_ ;
wire \sub3/insert_0/insert_2/_06_ ;
wire \sub3/insert_0/insert_2/_07_ ;
wire \sub3/insert_0/insert_3/_00_ ;
wire \sub3/insert_0/insert_3/_01_ ;
wire \sub3/insert_0/insert_3/_02_ ;
wire \sub3/insert_0/insert_3/_03_ ;
wire \sub3/insert_0/insert_3/_04_ ;
wire \sub3/insert_0/insert_3/_05_ ;
wire \sub3/insert_0/insert_3/_06_ ;
wire \sub3/insert_0/insert_3/_07_ ;
wire \xor3/_00_ ;
wire \xor3/_01_ ;
wire \xor3/_02_ ;
wire \xor3/_03_ ;
wire \xor3/_04_ ;
wire \xor3/_05_ ;
wire \xor3/_06_ ;
wire \xor3/_07_ ;
wire \xor3/_08_ ;
wire \xor3/_09_ ;
wire \xor3/_10_ ;
wire \xor3/_11_ ;
wire \xor3/_12_ ;
wire [2:0] BTN ;
wire [6:0] LD ;
wire [3:0] SW1 ;
wire [3:0] SW2 ;
wire [6:0] resul0 ;
wire [6:0] resul1 ;
wire [6:0] resul2 ;
wire [6:0] resul3 ;
wire [6:0] resul4 ;
wire [6:0] resul5 ;
wire [6:0] resul6 ;
wire [6:0] resul7 ;
wire [2:0] \sub3/SW0s ;


INV_X32 _134_ ( .A(_002_ ), .ZN(_047_ ) );
NOR2_X4 _135_ ( .A1(_047_ ), .A2(_001_ ), .ZN(_048_ ) );
AND3_X1 _136_ ( .A1(_048_ ), .A2(_000_ ), .A3(_113_ ), .ZN(_049_ ) );
INV_X2 _137_ ( .A(_000_ ), .ZN(_050_ ) );
AND2_X2 _138_ ( .A1(_048_ ), .A2(_050_ ), .ZN(_051_ ) );
AOI21_X1 _139_ ( .A(_049_ ), .B1(_106_ ), .B2(_051_ ), .ZN(_052_ ) );
INV_X32 _140_ ( .A(_001_ ), .ZN(_053_ ) );
NOR2_X4 _141_ ( .A1(_053_ ), .A2(_002_ ), .ZN(_054_ ) );
AND3_X1 _142_ ( .A1(_054_ ), .A2(_000_ ), .A3(_099_ ), .ZN(_055_ ) );
AND2_X2 _143_ ( .A1(_054_ ), .A2(_050_ ), .ZN(_056_ ) );
AOI21_X1 _144_ ( .A(_055_ ), .B1(_092_ ), .B2(_056_ ), .ZN(_057_ ) );
AND4_X1 _145_ ( .A1(_053_ ), .A2(_047_ ), .A3(_000_ ), .A4(_085_ ), .ZN(_058_ ) );
NOR2_X1 _146_ ( .A1(_001_ ), .A2(_002_ ), .ZN(_059_ ) );
AND2_X2 _147_ ( .A1(_059_ ), .A2(_050_ ), .ZN(_060_ ) );
AOI21_X1 _148_ ( .A(_058_ ), .B1(_078_ ), .B2(_060_ ), .ZN(_061_ ) );
AND2_X4 _149_ ( .A1(_001_ ), .A2(_002_ ), .ZN(_062_ ) );
AND3_X2 _150_ ( .A1(_062_ ), .A2(_000_ ), .A3(_127_ ), .ZN(_063_ ) );
AND2_X4 _151_ ( .A1(_062_ ), .A2(_050_ ), .ZN(_064_ ) );
AOI21_X2 _152_ ( .A(_063_ ), .B1(_120_ ), .B2(_064_ ), .ZN(_065_ ) );
NAND4_X1 _153_ ( .A1(_052_ ), .A2(_057_ ), .A3(_061_ ), .A4(_065_ ), .ZN(_003_ ) );
AND3_X1 _154_ ( .A1(_048_ ), .A2(_000_ ), .A3(_114_ ), .ZN(_066_ ) );
AOI21_X1 _155_ ( .A(_066_ ), .B1(_107_ ), .B2(_051_ ), .ZN(_067_ ) );
AND3_X1 _156_ ( .A1(_054_ ), .A2(_000_ ), .A3(_100_ ), .ZN(_068_ ) );
AOI21_X1 _157_ ( .A(_068_ ), .B1(_093_ ), .B2(_056_ ), .ZN(_069_ ) );
AND4_X1 _158_ ( .A1(_053_ ), .A2(_047_ ), .A3(_000_ ), .A4(_086_ ), .ZN(_070_ ) );
AOI21_X1 _159_ ( .A(_070_ ), .B1(_079_ ), .B2(_060_ ), .ZN(_071_ ) );
AND3_X2 _160_ ( .A1(_062_ ), .A2(_000_ ), .A3(_128_ ), .ZN(_072_ ) );
AOI21_X2 _161_ ( .A(_072_ ), .B1(_121_ ), .B2(_064_ ), .ZN(_073_ ) );
NAND4_X1 _162_ ( .A1(_067_ ), .A2(_069_ ), .A3(_071_ ), .A4(_073_ ), .ZN(_004_ ) );
AND3_X1 _163_ ( .A1(_048_ ), .A2(_000_ ), .A3(_115_ ), .ZN(_074_ ) );
AOI21_X1 _164_ ( .A(_074_ ), .B1(_108_ ), .B2(_051_ ), .ZN(_075_ ) );
AND3_X1 _165_ ( .A1(_054_ ), .A2(_000_ ), .A3(_101_ ), .ZN(_076_ ) );
AOI21_X1 _166_ ( .A(_076_ ), .B1(_094_ ), .B2(_056_ ), .ZN(_077_ ) );
AND4_X1 _167_ ( .A1(_053_ ), .A2(_047_ ), .A3(_000_ ), .A4(_087_ ), .ZN(_010_ ) );
AOI21_X1 _168_ ( .A(_010_ ), .B1(_080_ ), .B2(_060_ ), .ZN(_011_ ) );
AND3_X2 _169_ ( .A1(_062_ ), .A2(_000_ ), .A3(_129_ ), .ZN(_012_ ) );
AOI21_X2 _170_ ( .A(_012_ ), .B1(_122_ ), .B2(_064_ ), .ZN(_013_ ) );
NAND4_X1 _171_ ( .A1(_075_ ), .A2(_077_ ), .A3(_011_ ), .A4(_013_ ), .ZN(_005_ ) );
AND3_X1 _172_ ( .A1(_054_ ), .A2(_000_ ), .A3(_102_ ), .ZN(_014_ ) );
AOI21_X1 _173_ ( .A(_014_ ), .B1(_095_ ), .B2(_056_ ), .ZN(_015_ ) );
AND3_X2 _174_ ( .A1(_062_ ), .A2(_000_ ), .A3(_130_ ), .ZN(_016_ ) );
AOI21_X2 _175_ ( .A(_016_ ), .B1(_109_ ), .B2(_051_ ), .ZN(_017_ ) );
AND3_X2 _176_ ( .A1(_062_ ), .A2(_050_ ), .A3(_123_ ), .ZN(_018_ ) );
AND2_X1 _177_ ( .A1(_048_ ), .A2(_000_ ), .ZN(_019_ ) );
AOI21_X2 _178_ ( .A(_018_ ), .B1(_116_ ), .B2(_019_ ), .ZN(_020_ ) );
AND4_X1 _179_ ( .A1(_053_ ), .A2(_047_ ), .A3(_000_ ), .A4(_088_ ), .ZN(_021_ ) );
AOI21_X1 _180_ ( .A(_021_ ), .B1(_081_ ), .B2(_060_ ), .ZN(_022_ ) );
NAND4_X1 _181_ ( .A1(_015_ ), .A2(_017_ ), .A3(_020_ ), .A4(_022_ ), .ZN(_006_ ) );
AND3_X1 _182_ ( .A1(_048_ ), .A2(_050_ ), .A3(_110_ ), .ZN(_023_ ) );
AOI21_X1 _183_ ( .A(_023_ ), .B1(_117_ ), .B2(_019_ ), .ZN(_024_ ) );
AND3_X1 _184_ ( .A1(_054_ ), .A2(_000_ ), .A3(_103_ ), .ZN(_025_ ) );
AOI21_X1 _185_ ( .A(_025_ ), .B1(_096_ ), .B2(_056_ ), .ZN(_026_ ) );
AND4_X1 _186_ ( .A1(_053_ ), .A2(_047_ ), .A3(_000_ ), .A4(_089_ ), .ZN(_027_ ) );
AOI21_X1 _187_ ( .A(_027_ ), .B1(_082_ ), .B2(_060_ ), .ZN(_028_ ) );
AND3_X2 _188_ ( .A1(_062_ ), .A2(_000_ ), .A3(_131_ ), .ZN(_029_ ) );
AOI21_X2 _189_ ( .A(_029_ ), .B1(_124_ ), .B2(_064_ ), .ZN(_030_ ) );
NAND4_X1 _190_ ( .A1(_024_ ), .A2(_026_ ), .A3(_028_ ), .A4(_030_ ), .ZN(_007_ ) );
AND3_X1 _191_ ( .A1(_048_ ), .A2(_000_ ), .A3(_118_ ), .ZN(_031_ ) );
AOI21_X1 _192_ ( .A(_031_ ), .B1(_111_ ), .B2(_051_ ), .ZN(_032_ ) );
AND3_X1 _193_ ( .A1(_054_ ), .A2(_000_ ), .A3(_104_ ), .ZN(_033_ ) );
AOI21_X1 _194_ ( .A(_033_ ), .B1(_097_ ), .B2(_056_ ), .ZN(_034_ ) );
AND4_X1 _195_ ( .A1(_053_ ), .A2(_047_ ), .A3(_000_ ), .A4(_090_ ), .ZN(_035_ ) );
AOI21_X1 _196_ ( .A(_035_ ), .B1(_083_ ), .B2(_060_ ), .ZN(_036_ ) );
AND3_X2 _197_ ( .A1(_062_ ), .A2(_000_ ), .A3(_132_ ), .ZN(_037_ ) );
AOI21_X2 _198_ ( .A(_037_ ), .B1(_125_ ), .B2(_064_ ), .ZN(_038_ ) );
NAND4_X1 _199_ ( .A1(_032_ ), .A2(_034_ ), .A3(_036_ ), .A4(_038_ ), .ZN(_008_ ) );
AND3_X1 _200_ ( .A1(_048_ ), .A2(_000_ ), .A3(_119_ ), .ZN(_039_ ) );
AOI21_X1 _201_ ( .A(_039_ ), .B1(_112_ ), .B2(_051_ ), .ZN(_040_ ) );
AND3_X1 _202_ ( .A1(_054_ ), .A2(_000_ ), .A3(_105_ ), .ZN(_041_ ) );
AOI21_X1 _203_ ( .A(_041_ ), .B1(_098_ ), .B2(_056_ ), .ZN(_042_ ) );
AND4_X1 _204_ ( .A1(_053_ ), .A2(_047_ ), .A3(_000_ ), .A4(_091_ ), .ZN(_043_ ) );
AOI21_X1 _205_ ( .A(_043_ ), .B1(_084_ ), .B2(_060_ ), .ZN(_044_ ) );
AND3_X2 _206_ ( .A1(_062_ ), .A2(_000_ ), .A3(_133_ ), .ZN(_045_ ) );
AOI21_X2 _207_ ( .A(_045_ ), .B1(_126_ ), .B2(_064_ ), .ZN(_046_ ) );
NAND4_X1 _208_ ( .A1(_040_ ), .A2(_042_ ), .A3(_044_ ), .A4(_046_ ), .ZN(_009_ ) );
BUF_X1 _209_ ( .A(\BTN [1] ), .Z(_001_ ) );
BUF_X1 _210_ ( .A(\BTN [2] ), .Z(_002_ ) );
BUF_X1 _211_ ( .A(\BTN [0] ), .Z(_000_ ) );
BUF_X1 _212_ ( .A(\resul0 [0] ), .Z(_078_ ) );
BUF_X1 _213_ ( .A(\resul1 [0] ), .Z(_085_ ) );
BUF_X1 _214_ ( .A(\resul2 [0] ), .Z(_092_ ) );
BUF_X1 _215_ ( .A(\resul3 [0] ), .Z(_099_ ) );
BUF_X1 _216_ ( .A(\resul4 [0] ), .Z(_106_ ) );
BUF_X1 _217_ ( .A(\resul5 [0] ), .Z(_113_ ) );
BUF_X1 _218_ ( .A(\resul6 [0] ), .Z(_120_ ) );
BUF_X1 _219_ ( .A(\resul7 [0] ), .Z(_127_ ) );
BUF_X1 _220_ ( .A(_003_ ), .Z(\LD [0] ) );
BUF_X1 _221_ ( .A(\resul0 [1] ), .Z(_079_ ) );
BUF_X1 _222_ ( .A(\resul1 [1] ), .Z(_086_ ) );
BUF_X1 _223_ ( .A(\resul2 [1] ), .Z(_093_ ) );
BUF_X1 _224_ ( .A(\resul3 [1] ), .Z(_100_ ) );
BUF_X1 _225_ ( .A(\resul4 [1] ), .Z(_107_ ) );
BUF_X1 _226_ ( .A(\resul5 [1] ), .Z(_114_ ) );
BUF_X1 _227_ ( .A(\resul6 [1] ), .Z(_121_ ) );
BUF_X1 _228_ ( .A(\resul7 [1] ), .Z(_128_ ) );
BUF_X1 _229_ ( .A(_004_ ), .Z(\LD [1] ) );
BUF_X1 _230_ ( .A(\resul0 [2] ), .Z(_080_ ) );
BUF_X1 _231_ ( .A(\resul1 [2] ), .Z(_087_ ) );
BUF_X1 _232_ ( .A(\resul2 [2] ), .Z(_094_ ) );
BUF_X1 _233_ ( .A(\resul3 [2] ), .Z(_101_ ) );
BUF_X1 _234_ ( .A(\resul4 [2] ), .Z(_108_ ) );
BUF_X1 _235_ ( .A(\resul5 [2] ), .Z(_115_ ) );
BUF_X1 _236_ ( .A(\resul6 [2] ), .Z(_122_ ) );
BUF_X1 _237_ ( .A(\resul7 [2] ), .Z(_129_ ) );
BUF_X1 _238_ ( .A(_005_ ), .Z(\LD [2] ) );
BUF_X1 _239_ ( .A(\resul0 [3] ), .Z(_081_ ) );
BUF_X1 _240_ ( .A(\resul1 [3] ), .Z(_088_ ) );
BUF_X1 _241_ ( .A(\resul2 [3] ), .Z(_095_ ) );
BUF_X1 _242_ ( .A(\resul3 [3] ), .Z(_102_ ) );
BUF_X1 _243_ ( .A(\resul4 [3] ), .Z(_109_ ) );
BUF_X1 _244_ ( .A(\resul5 [3] ), .Z(_116_ ) );
BUF_X1 _245_ ( .A(\resul6 [3] ), .Z(_123_ ) );
BUF_X1 _246_ ( .A(\resul7 [3] ), .Z(_130_ ) );
BUF_X1 _247_ ( .A(_006_ ), .Z(\LD [3] ) );
BUF_X1 _248_ ( .A(\resul0 [4] ), .Z(_082_ ) );
BUF_X1 _249_ ( .A(\resul1 [4] ), .Z(_089_ ) );
BUF_X1 _250_ ( .A(\resul2 [4] ), .Z(_096_ ) );
BUF_X1 _251_ ( .A(\resul3 [4] ), .Z(_103_ ) );
BUF_X1 _252_ ( .A(\resul4 [4] ), .Z(_110_ ) );
BUF_X1 _253_ ( .A(\resul5 [4] ), .Z(_117_ ) );
BUF_X1 _254_ ( .A(\resul6 [4] ), .Z(_124_ ) );
BUF_X1 _255_ ( .A(\resul7 [4] ), .Z(_131_ ) );
BUF_X1 _256_ ( .A(_007_ ), .Z(\LD [4] ) );
BUF_X1 _257_ ( .A(\resul0 [5] ), .Z(_083_ ) );
BUF_X1 _258_ ( .A(\resul1 [5] ), .Z(_090_ ) );
BUF_X1 _259_ ( .A(\resul2 [5] ), .Z(_097_ ) );
BUF_X1 _260_ ( .A(\resul3 [5] ), .Z(_104_ ) );
BUF_X1 _261_ ( .A(\resul4 [5] ), .Z(_111_ ) );
BUF_X1 _262_ ( .A(\resul5 [5] ), .Z(_118_ ) );
BUF_X1 _263_ ( .A(\resul6 [5] ), .Z(_125_ ) );
BUF_X1 _264_ ( .A(\resul7 [5] ), .Z(_132_ ) );
BUF_X1 _265_ ( .A(_008_ ), .Z(\LD [5] ) );
BUF_X1 _266_ ( .A(\resul0 [6] ), .Z(_084_ ) );
BUF_X1 _267_ ( .A(\resul1 [6] ), .Z(_091_ ) );
BUF_X1 _268_ ( .A(\resul2 [6] ), .Z(_098_ ) );
BUF_X1 _269_ ( .A(\resul3 [6] ), .Z(_105_ ) );
BUF_X1 _270_ ( .A(\resul4 [6] ), .Z(_112_ ) );
BUF_X1 _271_ ( .A(\resul5 [6] ), .Z(_119_ ) );
BUF_X1 _272_ ( .A(\resul6 [6] ), .Z(_126_ ) );
BUF_X1 _273_ ( .A(\resul7 [6] ), .Z(_133_ ) );
BUF_X1 _274_ ( .A(_009_ ), .Z(\LD [6] ) );
NOR3_X1 \add3/_08_ ( .A1(\add3/_05_ ), .A2(\add3/_04_ ), .A3(\add3/_06_ ), .ZN(\add3/_01_ ) );
XOR2_X1 \add3/_09_ ( .A(\add3/_03_ ), .B(\add3/_02_ ), .Z(\add3/_00_ ) );
LOGIC0_X1 \add3/_10_ ( .Z(\add3/_07_ ) );
BUF_X1 \add3/_11_ ( .A(\add3/s0 ), .Z(\resul0 [0] ) );
BUF_X1 \add3/_12_ ( .A(\add3/s1 ), .Z(\resul0 [1] ) );
BUF_X1 \add3/_13_ ( .A(\add3/s2 ), .Z(\resul0 [2] ) );
BUF_X1 \add3/_14_ ( .A(\add3/s3 ), .Z(\resul0 [3] ) );
BUF_X1 \add3/_15_ ( .A(\add3/cout4 ), .Z(\resul0 [4] ) );
BUF_X1 \add3/_16_ ( .A(\add3/s1 ), .Z(\add3/_05_ ) );
BUF_X1 \add3/_17_ ( .A(\add3/s0 ), .Z(\add3/_04_ ) );
BUF_X1 \add3/_18_ ( .A(\add3/s2 ), .Z(\add3/_06_ ) );
BUF_X1 \add3/_19_ ( .A(\add3/_01_ ), .Z(\resul0 [6] ) );
BUF_X1 \add3/_20_ ( .A(\add3/cout4 ), .Z(\add3/_03_ ) );
BUF_X1 \add3/_21_ ( .A(\add3/cout3 ), .Z(\add3/_02_ ) );
BUF_X1 \add3/_22_ ( .A(\add3/_00_ ), .Z(\resul0 [5] ) );
XOR2_X2 \add3/insert_0/_08_ ( .A(\add3/insert_0/_02_ ), .B(\add3/insert_0/_00_ ), .Z(\add3/insert_0/_04_ ) );
XOR2_X1 \add3/insert_0/_09_ ( .A(\add3/insert_0/_04_ ), .B(\add3/insert_0/_01_ ), .Z(\add3/insert_0/_07_ ) );
NAND2_X1 \add3/insert_0/_10_ ( .A1(\add3/insert_0/_04_ ), .A2(\add3/insert_0/_01_ ), .ZN(\add3/insert_0/_05_ ) );
NAND2_X1 \add3/insert_0/_11_ ( .A1(\add3/insert_0/_02_ ), .A2(\add3/insert_0/_00_ ), .ZN(\add3/insert_0/_06_ ) );
NAND2_X1 \add3/insert_0/_12_ ( .A1(\add3/insert_0/_05_ ), .A2(\add3/insert_0/_06_ ), .ZN(\add3/insert_0/_03_ ) );
BUF_X1 \add3/insert_0/_13_ ( .A(\add3/_07_ ), .Z(\add3/insert_0/_02_ ) );
BUF_X1 \add3/insert_0/_14_ ( .A(\SW1 [0] ), .Z(\add3/insert_0/_00_ ) );
BUF_X1 \add3/insert_0/_15_ ( .A(\SW2 [0] ), .Z(\add3/insert_0/_01_ ) );
BUF_X1 \add3/insert_0/_16_ ( .A(\add3/insert_0/_07_ ), .Z(\add3/s0 ) );
BUF_X1 \add3/insert_0/_17_ ( .A(\add3/insert_0/_03_ ), .Z(\add3/cout1 ) );
XOR2_X2 \add3/insert_1/_08_ ( .A(\add3/insert_1/_02_ ), .B(\add3/insert_1/_00_ ), .Z(\add3/insert_1/_04_ ) );
XOR2_X1 \add3/insert_1/_09_ ( .A(\add3/insert_1/_04_ ), .B(\add3/insert_1/_01_ ), .Z(\add3/insert_1/_07_ ) );
NAND2_X1 \add3/insert_1/_10_ ( .A1(\add3/insert_1/_04_ ), .A2(\add3/insert_1/_01_ ), .ZN(\add3/insert_1/_05_ ) );
NAND2_X1 \add3/insert_1/_11_ ( .A1(\add3/insert_1/_02_ ), .A2(\add3/insert_1/_00_ ), .ZN(\add3/insert_1/_06_ ) );
NAND2_X1 \add3/insert_1/_12_ ( .A1(\add3/insert_1/_05_ ), .A2(\add3/insert_1/_06_ ), .ZN(\add3/insert_1/_03_ ) );
BUF_X1 \add3/insert_1/_13_ ( .A(\add3/cout1 ), .Z(\add3/insert_1/_02_ ) );
BUF_X1 \add3/insert_1/_14_ ( .A(\SW1 [1] ), .Z(\add3/insert_1/_00_ ) );
BUF_X1 \add3/insert_1/_15_ ( .A(\SW2 [1] ), .Z(\add3/insert_1/_01_ ) );
BUF_X1 \add3/insert_1/_16_ ( .A(\add3/insert_1/_07_ ), .Z(\add3/s1 ) );
BUF_X1 \add3/insert_1/_17_ ( .A(\add3/insert_1/_03_ ), .Z(\add3/cout2 ) );
XOR2_X2 \add3/insert_2/_08_ ( .A(\add3/insert_2/_02_ ), .B(\add3/insert_2/_00_ ), .Z(\add3/insert_2/_04_ ) );
XOR2_X1 \add3/insert_2/_09_ ( .A(\add3/insert_2/_04_ ), .B(\add3/insert_2/_01_ ), .Z(\add3/insert_2/_07_ ) );
NAND2_X1 \add3/insert_2/_10_ ( .A1(\add3/insert_2/_04_ ), .A2(\add3/insert_2/_01_ ), .ZN(\add3/insert_2/_05_ ) );
NAND2_X1 \add3/insert_2/_11_ ( .A1(\add3/insert_2/_02_ ), .A2(\add3/insert_2/_00_ ), .ZN(\add3/insert_2/_06_ ) );
NAND2_X1 \add3/insert_2/_12_ ( .A1(\add3/insert_2/_05_ ), .A2(\add3/insert_2/_06_ ), .ZN(\add3/insert_2/_03_ ) );
BUF_X1 \add3/insert_2/_13_ ( .A(\add3/cout2 ), .Z(\add3/insert_2/_02_ ) );
BUF_X1 \add3/insert_2/_14_ ( .A(\SW1 [2] ), .Z(\add3/insert_2/_00_ ) );
BUF_X1 \add3/insert_2/_15_ ( .A(\SW2 [2] ), .Z(\add3/insert_2/_01_ ) );
BUF_X1 \add3/insert_2/_16_ ( .A(\add3/insert_2/_07_ ), .Z(\add3/s2 ) );
BUF_X1 \add3/insert_2/_17_ ( .A(\add3/insert_2/_03_ ), .Z(\add3/cout3 ) );
XOR2_X2 \add3/insert_3/_08_ ( .A(\add3/insert_3/_02_ ), .B(\add3/insert_3/_00_ ), .Z(\add3/insert_3/_04_ ) );
XOR2_X1 \add3/insert_3/_09_ ( .A(\add3/insert_3/_04_ ), .B(\add3/insert_3/_01_ ), .Z(\add3/insert_3/_07_ ) );
NAND2_X1 \add3/insert_3/_10_ ( .A1(\add3/insert_3/_04_ ), .A2(\add3/insert_3/_01_ ), .ZN(\add3/insert_3/_05_ ) );
NAND2_X1 \add3/insert_3/_11_ ( .A1(\add3/insert_3/_02_ ), .A2(\add3/insert_3/_00_ ), .ZN(\add3/insert_3/_06_ ) );
NAND2_X1 \add3/insert_3/_12_ ( .A1(\add3/insert_3/_05_ ), .A2(\add3/insert_3/_06_ ), .ZN(\add3/insert_3/_03_ ) );
BUF_X1 \add3/insert_3/_13_ ( .A(\add3/cout3 ), .Z(\add3/insert_3/_02_ ) );
BUF_X1 \add3/insert_3/_14_ ( .A(\SW1 [3] ), .Z(\add3/insert_3/_00_ ) );
BUF_X1 \add3/insert_3/_15_ ( .A(\SW2 [3] ), .Z(\add3/insert_3/_01_ ) );
BUF_X1 \add3/insert_3/_16_ ( .A(\add3/insert_3/_07_ ), .Z(\add3/s3 ) );
BUF_X1 \add3/insert_3/_17_ ( .A(\add3/insert_3/_03_ ), .Z(\add3/cout4 ) );
AND2_X4 \and3/_13_ ( .A1(\and3/_04_ ), .A2(\and3/_00_ ), .ZN(\and3/_08_ ) );
AND2_X4 \and3/_14_ ( .A1(\and3/_05_ ), .A2(\and3/_01_ ), .ZN(\and3/_09_ ) );
AND2_X4 \and3/_15_ ( .A1(\and3/_06_ ), .A2(\and3/_02_ ), .ZN(\and3/_10_ ) );
AND2_X4 \and3/_16_ ( .A1(\and3/_07_ ), .A2(\and3/_03_ ), .ZN(\and3/_11_ ) );
LOGIC0_X1 \and3/_17_ ( .Z(\and3/_12_ ) );
BUF_X1 \and3/_18_ ( .A(\and3/_12_ ), .Z(\resul3 [4] ) );
BUF_X1 \and3/_19_ ( .A(\and3/_12_ ), .Z(\resul3 [5] ) );
BUF_X1 \and3/_20_ ( .A(\and3/_12_ ), .Z(\resul3 [6] ) );
BUF_X1 \and3/_21_ ( .A(\SW2 [0] ), .Z(\and3/_04_ ) );
BUF_X1 \and3/_22_ ( .A(\SW1 [0] ), .Z(\and3/_00_ ) );
BUF_X1 \and3/_23_ ( .A(\and3/_08_ ), .Z(\resul3 [0] ) );
BUF_X1 \and3/_24_ ( .A(\SW2 [1] ), .Z(\and3/_05_ ) );
BUF_X1 \and3/_25_ ( .A(\SW1 [1] ), .Z(\and3/_01_ ) );
BUF_X1 \and3/_26_ ( .A(\and3/_09_ ), .Z(\resul3 [1] ) );
BUF_X1 \and3/_27_ ( .A(\SW2 [2] ), .Z(\and3/_06_ ) );
BUF_X1 \and3/_28_ ( .A(\SW1 [2] ), .Z(\and3/_02_ ) );
BUF_X1 \and3/_29_ ( .A(\and3/_10_ ), .Z(\resul3 [2] ) );
BUF_X1 \and3/_30_ ( .A(\SW2 [3] ), .Z(\and3/_07_ ) );
BUF_X1 \and3/_31_ ( .A(\SW1 [3] ), .Z(\and3/_03_ ) );
BUF_X1 \and3/_32_ ( .A(\and3/_11_ ), .Z(\resul3 [3] ) );
INV_X32 \c3/_22_ ( .A(\c3/_04_ ), .ZN(\c3/_09_ ) );
AND2_X4 \c3/_23_ ( .A1(\c3/_09_ ), .A2(\c3/_07_ ), .ZN(\c3/_10_ ) );
INV_X32 \c3/_24_ ( .A(\c3/_03_ ), .ZN(\c3/_11_ ) );
AOI21_X4 \c3/_25_ ( .A(\c3/_10_ ), .B1(\c3/_11_ ), .B2(\c3/_06_ ), .ZN(\c3/_12_ ) );
NOR2_X1 \c3/_26_ ( .A1(\c3/_09_ ), .A2(\c3/_07_ ), .ZN(\c3/_13_ ) );
NOR2_X1 \c3/_27_ ( .A1(\c3/_11_ ), .A2(\c3/_06_ ), .ZN(\c3/_14_ ) );
NOR2_X1 \c3/_28_ ( .A1(\c3/_13_ ), .A2(\c3/_14_ ), .ZN(\c3/_15_ ) );
INV_X1 \c3/_29_ ( .A(\c3/_02_ ), .ZN(\c3/_16_ ) );
NOR2_X1 \c3/_30_ ( .A1(\c3/_16_ ), .A2(\c3/_05_ ), .ZN(\c3/_17_ ) );
INV_X1 \c3/_31_ ( .A(\c3/_17_ ), .ZN(\c3/_18_ ) );
AND2_X1 \c3/_32_ ( .A1(\c3/_16_ ), .A2(\c3/_05_ ), .ZN(\c3/_19_ ) );
INV_X1 \c3/_33_ ( .A(\c3/_19_ ), .ZN(\c3/_20_ ) );
AND4_X2 \c3/_34_ ( .A1(\c3/_12_ ), .A2(\c3/_15_ ), .A3(\c3/_18_ ), .A4(\c3/_20_ ), .ZN(\c3/_08_ ) );
NAND2_X1 \c3/_35_ ( .A1(\c3/_12_ ), .A2(\c3/_15_ ), .ZN(\c3/_21_ ) );
OAI22_X1 \c3/_36_ ( .A1(\c3/_21_ ), .A2(\c3/_18_ ), .B1(\c3/_10_ ), .B2(\c3/_15_ ), .ZN(\c3/_01_ ) );
OAI22_X1 \c3/_37_ ( .A1(\c3/_21_ ), .A2(\c3/_20_ ), .B1(\c3/_12_ ), .B2(\c3/_13_ ), .ZN(\c3/_00_ ) );
BUF_X1 \c3/_38_ ( .A(\resul6 [2] ), .Z(\resul6 [0] ) );
BUF_X1 \c3/_39_ ( .A(\resul6 [2] ), .Z(\resul6 [1] ) );
BUF_X1 \c3/_40_ ( .A(\c3/eq0 ), .Z(\resul6 [3] ) );
BUF_X1 \c3/_41_ ( .A(\resul6 [6] ), .Z(\resul6 [4] ) );
BUF_X1 \c3/_42_ ( .A(\resul6 [6] ), .Z(\resul6 [5] ) );
BUF_X1 \c3/_43_ ( .A(\SW1 [2] ), .Z(\c3/_04_ ) );
BUF_X1 \c3/_44_ ( .A(\SW2 [2] ), .Z(\c3/_07_ ) );
BUF_X1 \c3/_45_ ( .A(\SW1 [1] ), .Z(\c3/_03_ ) );
BUF_X1 \c3/_46_ ( .A(\SW2 [1] ), .Z(\c3/_06_ ) );
BUF_X1 \c3/_47_ ( .A(\SW1 [0] ), .Z(\c3/_02_ ) );
BUF_X1 \c3/_48_ ( .A(\SW2 [0] ), .Z(\c3/_05_ ) );
BUF_X1 \c3/_49_ ( .A(\c3/_08_ ), .Z(\c3/eq0 ) );
BUF_X1 \c3/_50_ ( .A(\c3/_01_ ), .Z(\resul6 [6] ) );
BUF_X1 \c3/_51_ ( .A(\c3/_00_ ), .Z(\resul6 [2] ) );
XNOR2_X2 \eq3/_10_ ( .A(\eq3/_04_ ), .B(\eq3/_01_ ), .ZN(\eq3/_08_ ) );
XNOR2_X2 \eq3/_11_ ( .A(\eq3/_03_ ), .B(\eq3/_00_ ), .ZN(\eq3/_09_ ) );
XNOR2_X2 \eq3/_12_ ( .A(\eq3/_05_ ), .B(\eq3/_02_ ), .ZN(\eq3/_07_ ) );
AND3_X1 \eq3/_13_ ( .A1(\eq3/_08_ ), .A2(\eq3/_09_ ), .A3(\eq3/_07_ ), .ZN(\eq3/_06_ ) );
BUF_X1 \eq3/_14_ ( .A(\eq3/eq0 ), .Z(\resul7 [0] ) );
BUF_X1 \eq3/_15_ ( .A(\eq3/eq0 ), .Z(\resul7 [1] ) );
BUF_X1 \eq3/_16_ ( .A(\eq3/eq0 ), .Z(\resul7 [2] ) );
BUF_X1 \eq3/_17_ ( .A(\eq3/eq0 ), .Z(\resul7 [3] ) );
BUF_X1 \eq3/_18_ ( .A(\eq3/eq0 ), .Z(\resul7 [4] ) );
BUF_X1 \eq3/_19_ ( .A(\eq3/eq0 ), .Z(\resul7 [5] ) );
BUF_X1 \eq3/_20_ ( .A(\eq3/eq0 ), .Z(\resul7 [6] ) );
BUF_X1 \eq3/_21_ ( .A(\SW2 [2] ), .Z(\eq3/_05_ ) );
BUF_X1 \eq3/_22_ ( .A(\SW1 [2] ), .Z(\eq3/_02_ ) );
BUF_X1 \eq3/_23_ ( .A(\SW2 [1] ), .Z(\eq3/_04_ ) );
BUF_X1 \eq3/_24_ ( .A(\SW1 [1] ), .Z(\eq3/_01_ ) );
BUF_X1 \eq3/_25_ ( .A(\SW2 [0] ), .Z(\eq3/_03_ ) );
BUF_X1 \eq3/_26_ ( .A(\SW1 [0] ), .Z(\eq3/_00_ ) );
BUF_X1 \eq3/_27_ ( .A(\eq3/_06_ ), .Z(\eq3/eq0 ) );
INV_X1 \not3/_09_ ( .A(\not3/_00_ ), .ZN(\not3/_04_ ) );
INV_X1 \not3/_10_ ( .A(\not3/_01_ ), .ZN(\not3/_05_ ) );
INV_X1 \not3/_11_ ( .A(\not3/_02_ ), .ZN(\not3/_06_ ) );
INV_X1 \not3/_12_ ( .A(\not3/_03_ ), .ZN(\not3/_07_ ) );
LOGIC0_X1 \not3/_13_ ( .Z(\not3/_08_ ) );
BUF_X1 \not3/_14_ ( .A(\not3/_08_ ), .Z(\resul2 [4] ) );
BUF_X1 \not3/_15_ ( .A(\not3/_08_ ), .Z(\resul2 [5] ) );
BUF_X1 \not3/_16_ ( .A(\not3/_08_ ), .Z(\resul2 [6] ) );
BUF_X1 \not3/_17_ ( .A(\SW1 [0] ), .Z(\not3/_00_ ) );
BUF_X1 \not3/_18_ ( .A(\not3/_04_ ), .Z(\resul2 [0] ) );
BUF_X1 \not3/_19_ ( .A(\SW1 [1] ), .Z(\not3/_01_ ) );
BUF_X1 \not3/_20_ ( .A(\not3/_05_ ), .Z(\resul2 [1] ) );
BUF_X1 \not3/_21_ ( .A(\SW1 [2] ), .Z(\not3/_02_ ) );
BUF_X1 \not3/_22_ ( .A(\not3/_06_ ), .Z(\resul2 [2] ) );
BUF_X1 \not3/_23_ ( .A(\SW1 [3] ), .Z(\not3/_03_ ) );
BUF_X1 \not3/_24_ ( .A(\not3/_07_ ), .Z(\resul2 [3] ) );
OR2_X4 \or3/_13_ ( .A1(\or3/_04_ ), .A2(\or3/_00_ ), .ZN(\or3/_08_ ) );
OR2_X4 \or3/_14_ ( .A1(\or3/_05_ ), .A2(\or3/_01_ ), .ZN(\or3/_09_ ) );
OR2_X4 \or3/_15_ ( .A1(\or3/_06_ ), .A2(\or3/_02_ ), .ZN(\or3/_10_ ) );
OR2_X4 \or3/_16_ ( .A1(\or3/_07_ ), .A2(\or3/_03_ ), .ZN(\or3/_11_ ) );
LOGIC0_X1 \or3/_17_ ( .Z(\or3/_12_ ) );
BUF_X1 \or3/_18_ ( .A(\or3/_12_ ), .Z(\resul4 [4] ) );
BUF_X1 \or3/_19_ ( .A(\or3/_12_ ), .Z(\resul4 [5] ) );
BUF_X1 \or3/_20_ ( .A(\or3/_12_ ), .Z(\resul4 [6] ) );
BUF_X1 \or3/_21_ ( .A(\SW2 [0] ), .Z(\or3/_04_ ) );
BUF_X1 \or3/_22_ ( .A(\SW1 [0] ), .Z(\or3/_00_ ) );
BUF_X1 \or3/_23_ ( .A(\or3/_08_ ), .Z(\resul4 [0] ) );
BUF_X1 \or3/_24_ ( .A(\SW2 [1] ), .Z(\or3/_05_ ) );
BUF_X1 \or3/_25_ ( .A(\SW1 [1] ), .Z(\or3/_01_ ) );
BUF_X1 \or3/_26_ ( .A(\or3/_09_ ), .Z(\resul4 [1] ) );
BUF_X1 \or3/_27_ ( .A(\SW2 [2] ), .Z(\or3/_06_ ) );
BUF_X1 \or3/_28_ ( .A(\SW1 [2] ), .Z(\or3/_02_ ) );
BUF_X1 \or3/_29_ ( .A(\or3/_10_ ), .Z(\resul4 [2] ) );
BUF_X1 \or3/_30_ ( .A(\SW2 [3] ), .Z(\or3/_07_ ) );
BUF_X1 \or3/_31_ ( .A(\SW1 [3] ), .Z(\or3/_03_ ) );
BUF_X1 \or3/_32_ ( .A(\or3/_11_ ), .Z(\resul4 [3] ) );
XOR2_X1 \sub3/_07_ ( .A(\sub3/_03_ ), .B(\sub3/_02_ ), .Z(\sub3/_00_ ) );
NOR2_X4 \sub3/_08_ ( .A1(\sub3/_03_ ), .A2(\sub3/_02_ ), .ZN(\sub3/_05_ ) );
XNOR2_X1 \sub3/_09_ ( .A(\sub3/_05_ ), .B(\sub3/_04_ ), .ZN(\sub3/_01_ ) );
LOGIC1_X1 \sub3/_10_ ( .Z(\sub3/_06_ ) );
BUF_X1 \sub3/_11_ ( .A(\SW2 [0] ), .Z(\sub3/SW0s [0] ) );
BUF_X1 \sub3/_12_ ( .A(\SW2 [1] ), .Z(\sub3/_03_ ) );
BUF_X1 \sub3/_13_ ( .A(\SW2 [0] ), .Z(\sub3/_02_ ) );
BUF_X1 \sub3/_14_ ( .A(\sub3/_00_ ), .Z(\sub3/SW0s [1] ) );
BUF_X1 \sub3/_15_ ( .A(\SW2 [2] ), .Z(\sub3/_04_ ) );
BUF_X1 \sub3/_16_ ( .A(\sub3/_01_ ), .Z(\sub3/SW0s [2] ) );
NOR3_X1 \sub3/insert_0/_08_ ( .A1(\sub3/insert_0/_05_ ), .A2(\sub3/insert_0/_04_ ), .A3(\sub3/insert_0/_06_ ), .ZN(\sub3/insert_0/_01_ ) );
XOR2_X1 \sub3/insert_0/_09_ ( .A(\sub3/insert_0/_03_ ), .B(\sub3/insert_0/_02_ ), .Z(\sub3/insert_0/_00_ ) );
LOGIC0_X1 \sub3/insert_0/_10_ ( .Z(\sub3/insert_0/_07_ ) );
BUF_X1 \sub3/insert_0/_11_ ( .A(\sub3/insert_0/s0 ), .Z(\resul1 [0] ) );
BUF_X1 \sub3/insert_0/_12_ ( .A(\sub3/insert_0/s1 ), .Z(\resul1 [1] ) );
BUF_X1 \sub3/insert_0/_13_ ( .A(\sub3/insert_0/s2 ), .Z(\resul1 [2] ) );
BUF_X1 \sub3/insert_0/_14_ ( .A(\sub3/insert_0/s3 ), .Z(\resul1 [3] ) );
BUF_X1 \sub3/insert_0/_15_ ( .A(\sub3/insert_0/cout4 ), .Z(\resul1 [4] ) );
BUF_X1 \sub3/insert_0/_16_ ( .A(\sub3/insert_0/s1 ), .Z(\sub3/insert_0/_05_ ) );
BUF_X1 \sub3/insert_0/_17_ ( .A(\sub3/insert_0/s0 ), .Z(\sub3/insert_0/_04_ ) );
BUF_X1 \sub3/insert_0/_18_ ( .A(\sub3/insert_0/s2 ), .Z(\sub3/insert_0/_06_ ) );
BUF_X1 \sub3/insert_0/_19_ ( .A(\sub3/insert_0/_01_ ), .Z(\resul1 [6] ) );
BUF_X1 \sub3/insert_0/_20_ ( .A(\sub3/insert_0/cout4 ), .Z(\sub3/insert_0/_03_ ) );
BUF_X1 \sub3/insert_0/_21_ ( .A(\sub3/insert_0/cout3 ), .Z(\sub3/insert_0/_02_ ) );
BUF_X1 \sub3/insert_0/_22_ ( .A(\sub3/insert_0/_00_ ), .Z(\resul1 [5] ) );
XOR2_X2 \sub3/insert_0/insert_0/_08_ ( .A(\sub3/insert_0/insert_0/_02_ ), .B(\sub3/insert_0/insert_0/_00_ ), .Z(\sub3/insert_0/insert_0/_04_ ) );
XOR2_X1 \sub3/insert_0/insert_0/_09_ ( .A(\sub3/insert_0/insert_0/_04_ ), .B(\sub3/insert_0/insert_0/_01_ ), .Z(\sub3/insert_0/insert_0/_07_ ) );
NAND2_X1 \sub3/insert_0/insert_0/_10_ ( .A1(\sub3/insert_0/insert_0/_04_ ), .A2(\sub3/insert_0/insert_0/_01_ ), .ZN(\sub3/insert_0/insert_0/_05_ ) );
NAND2_X1 \sub3/insert_0/insert_0/_11_ ( .A1(\sub3/insert_0/insert_0/_02_ ), .A2(\sub3/insert_0/insert_0/_00_ ), .ZN(\sub3/insert_0/insert_0/_06_ ) );
NAND2_X1 \sub3/insert_0/insert_0/_12_ ( .A1(\sub3/insert_0/insert_0/_05_ ), .A2(\sub3/insert_0/insert_0/_06_ ), .ZN(\sub3/insert_0/insert_0/_03_ ) );
BUF_X1 \sub3/insert_0/insert_0/_13_ ( .A(\sub3/insert_0/_07_ ), .Z(\sub3/insert_0/insert_0/_02_ ) );
BUF_X1 \sub3/insert_0/insert_0/_14_ ( .A(\SW1 [0] ), .Z(\sub3/insert_0/insert_0/_00_ ) );
BUF_X1 \sub3/insert_0/insert_0/_15_ ( .A(\SW2 [0] ), .Z(\sub3/insert_0/insert_0/_01_ ) );
BUF_X1 \sub3/insert_0/insert_0/_16_ ( .A(\sub3/insert_0/insert_0/_07_ ), .Z(\sub3/insert_0/s0 ) );
BUF_X1 \sub3/insert_0/insert_0/_17_ ( .A(\sub3/insert_0/insert_0/_03_ ), .Z(\sub3/insert_0/cout1 ) );
XOR2_X2 \sub3/insert_0/insert_1/_08_ ( .A(\sub3/insert_0/insert_1/_02_ ), .B(\sub3/insert_0/insert_1/_00_ ), .Z(\sub3/insert_0/insert_1/_04_ ) );
XOR2_X1 \sub3/insert_0/insert_1/_09_ ( .A(\sub3/insert_0/insert_1/_04_ ), .B(\sub3/insert_0/insert_1/_01_ ), .Z(\sub3/insert_0/insert_1/_07_ ) );
NAND2_X1 \sub3/insert_0/insert_1/_10_ ( .A1(\sub3/insert_0/insert_1/_04_ ), .A2(\sub3/insert_0/insert_1/_01_ ), .ZN(\sub3/insert_0/insert_1/_05_ ) );
NAND2_X1 \sub3/insert_0/insert_1/_11_ ( .A1(\sub3/insert_0/insert_1/_02_ ), .A2(\sub3/insert_0/insert_1/_00_ ), .ZN(\sub3/insert_0/insert_1/_06_ ) );
NAND2_X1 \sub3/insert_0/insert_1/_12_ ( .A1(\sub3/insert_0/insert_1/_05_ ), .A2(\sub3/insert_0/insert_1/_06_ ), .ZN(\sub3/insert_0/insert_1/_03_ ) );
BUF_X1 \sub3/insert_0/insert_1/_13_ ( .A(\sub3/insert_0/cout1 ), .Z(\sub3/insert_0/insert_1/_02_ ) );
BUF_X1 \sub3/insert_0/insert_1/_14_ ( .A(\SW1 [1] ), .Z(\sub3/insert_0/insert_1/_00_ ) );
BUF_X1 \sub3/insert_0/insert_1/_15_ ( .A(\sub3/SW0s [1] ), .Z(\sub3/insert_0/insert_1/_01_ ) );
BUF_X1 \sub3/insert_0/insert_1/_16_ ( .A(\sub3/insert_0/insert_1/_07_ ), .Z(\sub3/insert_0/s1 ) );
BUF_X1 \sub3/insert_0/insert_1/_17_ ( .A(\sub3/insert_0/insert_1/_03_ ), .Z(\sub3/insert_0/cout2 ) );
XOR2_X2 \sub3/insert_0/insert_2/_08_ ( .A(\sub3/insert_0/insert_2/_02_ ), .B(\sub3/insert_0/insert_2/_00_ ), .Z(\sub3/insert_0/insert_2/_04_ ) );
XOR2_X1 \sub3/insert_0/insert_2/_09_ ( .A(\sub3/insert_0/insert_2/_04_ ), .B(\sub3/insert_0/insert_2/_01_ ), .Z(\sub3/insert_0/insert_2/_07_ ) );
NAND2_X1 \sub3/insert_0/insert_2/_10_ ( .A1(\sub3/insert_0/insert_2/_04_ ), .A2(\sub3/insert_0/insert_2/_01_ ), .ZN(\sub3/insert_0/insert_2/_05_ ) );
NAND2_X1 \sub3/insert_0/insert_2/_11_ ( .A1(\sub3/insert_0/insert_2/_02_ ), .A2(\sub3/insert_0/insert_2/_00_ ), .ZN(\sub3/insert_0/insert_2/_06_ ) );
NAND2_X1 \sub3/insert_0/insert_2/_12_ ( .A1(\sub3/insert_0/insert_2/_05_ ), .A2(\sub3/insert_0/insert_2/_06_ ), .ZN(\sub3/insert_0/insert_2/_03_ ) );
BUF_X1 \sub3/insert_0/insert_2/_13_ ( .A(\sub3/insert_0/cout2 ), .Z(\sub3/insert_0/insert_2/_02_ ) );
BUF_X1 \sub3/insert_0/insert_2/_14_ ( .A(\SW1 [2] ), .Z(\sub3/insert_0/insert_2/_00_ ) );
BUF_X1 \sub3/insert_0/insert_2/_15_ ( .A(\sub3/SW0s [2] ), .Z(\sub3/insert_0/insert_2/_01_ ) );
BUF_X1 \sub3/insert_0/insert_2/_16_ ( .A(\sub3/insert_0/insert_2/_07_ ), .Z(\sub3/insert_0/s2 ) );
BUF_X1 \sub3/insert_0/insert_2/_17_ ( .A(\sub3/insert_0/insert_2/_03_ ), .Z(\sub3/insert_0/cout3 ) );
XOR2_X2 \sub3/insert_0/insert_3/_08_ ( .A(\sub3/insert_0/insert_3/_02_ ), .B(\sub3/insert_0/insert_3/_00_ ), .Z(\sub3/insert_0/insert_3/_04_ ) );
XOR2_X1 \sub3/insert_0/insert_3/_09_ ( .A(\sub3/insert_0/insert_3/_04_ ), .B(\sub3/insert_0/insert_3/_01_ ), .Z(\sub3/insert_0/insert_3/_07_ ) );
NAND2_X1 \sub3/insert_0/insert_3/_10_ ( .A1(\sub3/insert_0/insert_3/_04_ ), .A2(\sub3/insert_0/insert_3/_01_ ), .ZN(\sub3/insert_0/insert_3/_05_ ) );
NAND2_X1 \sub3/insert_0/insert_3/_11_ ( .A1(\sub3/insert_0/insert_3/_02_ ), .A2(\sub3/insert_0/insert_3/_00_ ), .ZN(\sub3/insert_0/insert_3/_06_ ) );
NAND2_X1 \sub3/insert_0/insert_3/_12_ ( .A1(\sub3/insert_0/insert_3/_05_ ), .A2(\sub3/insert_0/insert_3/_06_ ), .ZN(\sub3/insert_0/insert_3/_03_ ) );
BUF_X1 \sub3/insert_0/insert_3/_13_ ( .A(\sub3/insert_0/cout3 ), .Z(\sub3/insert_0/insert_3/_02_ ) );
BUF_X1 \sub3/insert_0/insert_3/_14_ ( .A(\SW1 [3] ), .Z(\sub3/insert_0/insert_3/_00_ ) );
BUF_X1 \sub3/insert_0/insert_3/_15_ ( .A(\sub3/_06_ ), .Z(\sub3/insert_0/insert_3/_01_ ) );
BUF_X1 \sub3/insert_0/insert_3/_16_ ( .A(\sub3/insert_0/insert_3/_07_ ), .Z(\sub3/insert_0/s3 ) );
BUF_X1 \sub3/insert_0/insert_3/_17_ ( .A(\sub3/insert_0/insert_3/_03_ ), .Z(\sub3/insert_0/cout4 ) );
XOR2_X1 \xor3/_13_ ( .A(\xor3/_04_ ), .B(\xor3/_00_ ), .Z(\xor3/_08_ ) );
XOR2_X1 \xor3/_14_ ( .A(\xor3/_05_ ), .B(\xor3/_01_ ), .Z(\xor3/_09_ ) );
XOR2_X1 \xor3/_15_ ( .A(\xor3/_06_ ), .B(\xor3/_02_ ), .Z(\xor3/_10_ ) );
XOR2_X1 \xor3/_16_ ( .A(\xor3/_07_ ), .B(\xor3/_03_ ), .Z(\xor3/_11_ ) );
LOGIC0_X1 \xor3/_17_ ( .Z(\xor3/_12_ ) );
BUF_X1 \xor3/_18_ ( .A(\xor3/_12_ ), .Z(\resul5 [4] ) );
BUF_X1 \xor3/_19_ ( .A(\xor3/_12_ ), .Z(\resul5 [5] ) );
BUF_X1 \xor3/_20_ ( .A(\xor3/_12_ ), .Z(\resul5 [6] ) );
BUF_X1 \xor3/_21_ ( .A(\SW2 [0] ), .Z(\xor3/_04_ ) );
BUF_X1 \xor3/_22_ ( .A(\SW1 [0] ), .Z(\xor3/_00_ ) );
BUF_X1 \xor3/_23_ ( .A(\xor3/_08_ ), .Z(\resul5 [0] ) );
BUF_X1 \xor3/_24_ ( .A(\SW2 [1] ), .Z(\xor3/_05_ ) );
BUF_X1 \xor3/_25_ ( .A(\SW1 [1] ), .Z(\xor3/_01_ ) );
BUF_X1 \xor3/_26_ ( .A(\xor3/_09_ ), .Z(\resul5 [1] ) );
BUF_X1 \xor3/_27_ ( .A(\SW2 [2] ), .Z(\xor3/_06_ ) );
BUF_X1 \xor3/_28_ ( .A(\SW1 [2] ), .Z(\xor3/_02_ ) );
BUF_X1 \xor3/_29_ ( .A(\xor3/_10_ ), .Z(\resul5 [2] ) );
BUF_X1 \xor3/_30_ ( .A(\SW2 [3] ), .Z(\xor3/_07_ ) );
BUF_X1 \xor3/_31_ ( .A(\SW1 [3] ), .Z(\xor3/_03_ ) );
BUF_X1 \xor3/_32_ ( .A(\xor3/_11_ ), .Z(\resul5 [3] ) );

endmodule
