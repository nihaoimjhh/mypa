//Generate the verilog at 2024-08-18T18:17:28
module top (
a,
s,
y
);

input [7:0] a ;
input [1:0] s ;
output [1:0] y ;

wire _0_ ;
wire _1_ ;
wire \i0/_0_ ;
wire \i0/i0/_00_ ;
wire \i0/i0/_01_ ;
wire \i0/i0/_02_ ;
wire \i0/i0/_03_ ;
wire \i0/i0/_04_ ;
wire \i0/i0/_05_ ;
wire \i0/i0/_06_ ;
wire \i0/i0/_07_ ;
wire \i0/i0/_08_ ;
wire \i0/i0/_09_ ;
wire \i0/i0/_10_ ;
wire \i0/i0/_11_ ;
wire \i0/i0/_12_ ;
wire \i0/i0/_13_ ;
wire \i0/i0/_14_ ;
wire \i0/i0/_15_ ;
wire \i0/i0/_16_ ;
wire \i0/i0/_17_ ;
wire \i0/i0/_18_ ;
wire \i0/i0/_19_ ;
wire \i0/i0/_20_ ;
wire \i0/i0/_21_ ;
wire \i0/i0/_22_ ;
wire \i0/i0/_23_ ;
wire \i0/i0/_24_ ;
wire \i0/i0/_25_ ;
wire \i0/i0/_26_ ;
wire \i0/i0/_27_ ;
wire \i0/i0/_28_ ;
wire \i0/i0/_29_ ;
wire \i0/i0/_30_ ;
wire \i0/i0/_31_ ;
wire \i0/i0/_32_ ;
wire \i0/i0/_33_ ;
wire \i0/i0/_34_ ;
wire \i0/i0/_35_ ;
wire \a[0] ;
wire \a[1] ;
wire \a[2] ;
wire \a[3] ;
wire \a[4] ;
wire \a[5] ;
wire \a[6] ;
wire \a[7] ;
wire \s[0] ;
wire \s[1] ;
wire \y[0] ;
wire \y[1] ;

assign \a[0] = a[0] ;
assign \a[1] = a[1] ;
assign \a[2] = a[2] ;
assign \a[3] = a[3] ;
assign \a[4] = a[4] ;
assign \a[5] = a[5] ;
assign \a[6] = a[6] ;
assign \a[7] = a[7] ;
assign \s[0] = s[0] ;
assign \s[1] = s[1] ;
assign y[0] = \y[0] ;
assign y[1] = \y[1] ;

LOGIC1_X1 _2_ ( .Z(_0_ ) );
LOGIC0_X1 _3_ ( .Z(_1_ ) );
LOGIC0_X1 \i0/_1_ ( .Z(\i0/_0_ ) );
XNOR2_X2 \i0/i0/_36_ ( .A(\i0/i0/_01_ ), .B(\i0/i0/_15_ ), .ZN(\i0/i0/_18_ ) );
XNOR2_X2 \i0/i0/_37_ ( .A(\i0/i0/_00_ ), .B(\i0/i0/_14_ ), .ZN(\i0/i0/_19_ ) );
NAND3_X1 \i0/i0/_38_ ( .A1(\i0/i0/_18_ ), .A2(\i0/i0/_19_ ), .A3(\i0/i0/_12_ ), .ZN(\i0/i0/_20_ ) );
XNOR2_X2 \i0/i0/_39_ ( .A(\i0/i0/_11_ ), .B(\i0/i0/_01_ ), .ZN(\i0/i0/_21_ ) );
XNOR2_X2 \i0/i0/_40_ ( .A(\i0/i0/_10_ ), .B(\i0/i0/_00_ ), .ZN(\i0/i0/_22_ ) );
NAND3_X1 \i0/i0/_41_ ( .A1(\i0/i0/_21_ ), .A2(\i0/i0/_22_ ), .A3(\i0/i0/_02_ ), .ZN(\i0/i0/_23_ ) );
XNOR2_X2 \i0/i0/_42_ ( .A(\i0/i0/_01_ ), .B(\i0/i0/_08_ ), .ZN(\i0/i0/_24_ ) );
XNOR2_X2 \i0/i0/_43_ ( .A(\i0/i0/_00_ ), .B(\i0/i0/_07_ ), .ZN(\i0/i0/_25_ ) );
NAND3_X1 \i0/i0/_44_ ( .A1(\i0/i0/_24_ ), .A2(\i0/i0/_25_ ), .A3(\i0/i0/_05_ ), .ZN(\i0/i0/_26_ ) );
XNOR2_X2 \i0/i0/_45_ ( .A(\i0/i0/_01_ ), .B(\i0/i0/_04_ ), .ZN(\i0/i0/_27_ ) );
XNOR2_X2 \i0/i0/_46_ ( .A(\i0/i0/_00_ ), .B(\i0/i0/_03_ ), .ZN(\i0/i0/_28_ ) );
NAND3_X1 \i0/i0/_47_ ( .A1(\i0/i0/_27_ ), .A2(\i0/i0/_28_ ), .A3(\i0/i0/_16_ ), .ZN(\i0/i0/_29_ ) );
NAND4_X1 \i0/i0/_48_ ( .A1(\i0/i0/_20_ ), .A2(\i0/i0/_23_ ), .A3(\i0/i0/_26_ ), .A4(\i0/i0/_29_ ), .ZN(\i0/i0/_34_ ) );
NAND3_X1 \i0/i0/_49_ ( .A1(\i0/i0/_18_ ), .A2(\i0/i0/_19_ ), .A3(\i0/i0/_13_ ), .ZN(\i0/i0/_30_ ) );
NAND3_X1 \i0/i0/_50_ ( .A1(\i0/i0/_21_ ), .A2(\i0/i0/_22_ ), .A3(\i0/i0/_09_ ), .ZN(\i0/i0/_31_ ) );
NAND3_X1 \i0/i0/_51_ ( .A1(\i0/i0/_24_ ), .A2(\i0/i0/_25_ ), .A3(\i0/i0/_06_ ), .ZN(\i0/i0/_32_ ) );
NAND3_X1 \i0/i0/_52_ ( .A1(\i0/i0/_27_ ), .A2(\i0/i0/_28_ ), .A3(\i0/i0/_17_ ), .ZN(\i0/i0/_33_ ) );
NAND4_X1 \i0/i0/_53_ ( .A1(\i0/i0/_30_ ), .A2(\i0/i0/_31_ ), .A3(\i0/i0/_32_ ), .A4(\i0/i0/_33_ ), .ZN(\i0/i0/_35_ ) );
BUF_X1 \i0/i0/_54_ ( .A(_0_ ), .Z(\i0/i0/_10_ ) );
BUF_X1 \i0/i0/_55_ ( .A(\s[0] ), .Z(\i0/i0/_00_ ) );
BUF_X1 \i0/i0/_56_ ( .A(_0_ ), .Z(\i0/i0/_11_ ) );
BUF_X1 \i0/i0/_57_ ( .A(\s[1] ), .Z(\i0/i0/_01_ ) );
BUF_X1 \i0/i0/_58_ ( .A(\a[6] ), .Z(\i0/i0/_02_ ) );
BUF_X1 \i0/i0/_59_ ( .A(_1_ ), .Z(\i0/i0/_14_ ) );
BUF_X1 \i0/i0/_60_ ( .A(_0_ ), .Z(\i0/i0/_15_ ) );
BUF_X1 \i0/i0/_61_ ( .A(\a[4] ), .Z(\i0/i0/_12_ ) );
BUF_X1 \i0/i0/_62_ ( .A(_0_ ), .Z(\i0/i0/_03_ ) );
BUF_X1 \i0/i0/_63_ ( .A(_1_ ), .Z(\i0/i0/_04_ ) );
BUF_X1 \i0/i0/_64_ ( .A(\a[2] ), .Z(\i0/i0/_16_ ) );
BUF_X1 \i0/i0/_65_ ( .A(_1_ ), .Z(\i0/i0/_07_ ) );
BUF_X1 \i0/i0/_66_ ( .A(_1_ ), .Z(\i0/i0/_08_ ) );
BUF_X1 \i0/i0/_67_ ( .A(\a[0] ), .Z(\i0/i0/_05_ ) );
BUF_X1 \i0/i0/_68_ ( .A(\i0/i0/_34_ ), .Z(\y[0] ) );
BUF_X1 \i0/i0/_69_ ( .A(\a[7] ), .Z(\i0/i0/_09_ ) );
BUF_X1 \i0/i0/_70_ ( .A(\a[5] ), .Z(\i0/i0/_13_ ) );
BUF_X1 \i0/i0/_71_ ( .A(\a[3] ), .Z(\i0/i0/_17_ ) );
BUF_X1 \i0/i0/_72_ ( .A(\a[1] ), .Z(\i0/i0/_06_ ) );
BUF_X1 \i0/i0/_73_ ( .A(\i0/i0/_35_ ), .Z(\y[1] ) );

endmodule
