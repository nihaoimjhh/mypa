//Generate the verilog at 2024-08-18T18:17:48
module top (
LD4,
LD,
SEG,
SEG0,
SW
);

output LD4 ;
output [2:0] LD ;
output [6:0] SEG ;
output [7:0] SEG0 ;
input [7:0] SW ;

wire _00_ ;
wire _01_ ;
wire _02_ ;
wire _03_ ;
wire _04_ ;
wire _05_ ;
wire _06_ ;
wire _07_ ;
wire _08_ ;
wire _09_ ;
wire _10_ ;
wire _11_ ;
wire _12_ ;
wire _13_ ;
wire _14_ ;
wire _15_ ;
wire _16_ ;
wire _17_ ;
wire _18_ ;
wire _19_ ;
wire _20_ ;
wire _21_ ;
wire _22_ ;
wire _23_ ;
wire _24_ ;
wire _25_ ;
wire _26_ ;
wire _27_ ;
wire _28_ ;
wire _29_ ;
wire _30_ ;
wire _31_ ;
wire _32_ ;
wire _33_ ;
wire LD4 ;
wire \LD[0] ;
wire \LD[1] ;
wire \LD[2] ;
wire \SEG[0] ;
wire \SEG[1] ;
wire \SEG[2] ;
wire \SEG[3] ;
wire \SEG[4] ;
wire \SEG[5] ;
wire \SEG[6] ;
wire \SEG0[0] ;
wire \SEG0[1] ;
wire \SEG0[2] ;
wire \SEG0[3] ;
wire \SEG0[4] ;
wire \SEG0[5] ;
wire \SEG0[6] ;
wire \SEG0[7] ;
wire \SW[0] ;
wire \SW[1] ;
wire \SW[2] ;
wire \SW[3] ;
wire \SW[4] ;
wire \SW[5] ;
wire \SW[6] ;
wire \SW[7] ;

assign LD[0] = \LD[0] ;
assign LD[1] = \LD[1] ;
assign LD[2] = \LD[2] ;
assign SEG[0] = \SEG[0] ;
assign SEG[1] = \SEG[1] ;
assign SEG[2] = \SEG[2] ;
assign SEG[3] = \SEG[3] ;
assign SEG[4] = \SEG[4] ;
assign SEG[5] = \SEG[5] ;
assign SEG[6] = \SEG[6] ;
assign SEG0[0] = \SEG0[0] ;
assign SEG0[1] = \SEG0[1] ;
assign SEG0[2] = \SEG0[2] ;
assign SEG0[3] = \SEG0[3] ;
assign SEG0[4] = \SEG0[4] ;
assign SEG0[5] = \SEG0[5] ;
assign SEG0[6] = \SEG0[6] ;
assign SEG0[7] = \SEG0[7] ;
assign \SW[1] = SW[1] ;
assign \SW[2] = SW[2] ;
assign \SW[3] = SW[3] ;
assign \SW[4] = SW[4] ;
assign \SW[5] = SW[5] ;
assign \SW[6] = SW[6] ;
assign \SW[7] = SW[7] ;

INV_X32 _34_ ( .A(_16_ ), .ZN(_18_ ) );
INV_X16 _35_ ( .A(_17_ ), .ZN(_19_ ) );
INV_X32 _36_ ( .A(_15_ ), .ZN(_20_ ) );
NAND3_X4 _37_ ( .A1(_18_ ), .A2(_19_ ), .A3(_20_ ), .ZN(_21_ ) );
NOR3_X4 _38_ ( .A1(_21_ ), .A2(_14_ ), .A3(_13_ ), .ZN(_22_ ) );
INV_X1 _39_ ( .A(_12_ ), .ZN(_23_ ) );
INV_X1 _40_ ( .A(_11_ ), .ZN(_24_ ) );
AND3_X1 _41_ ( .A1(_22_ ), .A2(_23_ ), .A3(_24_ ), .ZN(_25_ ) );
INV_X1 _42_ ( .A(_25_ ), .ZN(_00_ ) );
NOR2_X2 _43_ ( .A1(_21_ ), .A2(_14_ ), .ZN(_26_ ) );
INV_X1 _44_ ( .A(_26_ ), .ZN(_03_ ) );
AND2_X4 _45_ ( .A1(_22_ ), .A2(_12_ ), .ZN(_08_ ) );
AND2_X4 _46_ ( .A1(_26_ ), .A2(_13_ ), .ZN(_27_ ) );
OR4_X2 _47_ ( .A1(_16_ ), .A2(_08_ ), .A3(_17_ ), .A4(_27_ ), .ZN(_02_ ) );
AND3_X2 _48_ ( .A1(_22_ ), .A2(_23_ ), .A3(_11_ ), .ZN(_28_ ) );
NOR2_X1 _49_ ( .A1(_28_ ), .A2(_27_ ), .ZN(_29_ ) );
OAI211_X2 _50_ ( .A(_29_ ), .B(_19_ ), .C1(_16_ ), .C2(_20_ ), .ZN(_01_ ) );
AND2_X1 _51_ ( .A1(_22_ ), .A2(_23_ ), .ZN(_30_ ) );
AOI221_X1 _52_ ( .A(_08_ ), .B1(_16_ ), .B2(_19_ ), .C1(_24_ ), .C2(_30_ ), .ZN(_06_ ) );
INV_X1 _53_ ( .A(_28_ ), .ZN(_31_ ) );
NAND4_X1 _54_ ( .A1(_18_ ), .A2(_19_ ), .A3(_20_ ), .A4(_14_ ), .ZN(_32_ ) );
NAND2_X1 _55_ ( .A1(_31_ ), .A2(_32_ ), .ZN(_10_ ) );
AOI21_X1 _56_ ( .A(_17_ ), .B1(_18_ ), .B2(_20_ ), .ZN(_09_ ) );
NAND3_X1 _57_ ( .A1(_31_ ), .A2(_19_ ), .A3(_32_ ), .ZN(_07_ ) );
OR4_X2 _58_ ( .A1(_17_ ), .A2(_28_ ), .A3(_08_ ), .A4(_27_ ), .ZN(_05_ ) );
OR2_X1 _59_ ( .A1(_30_ ), .A2(_17_ ), .ZN(_04_ ) );
LOGIC1_X1 _60_ ( .Z(_33_ ) );
BUF_X1 _61_ ( .A(_33_ ), .Z(\SEG0[0] ) );
BUF_X1 _62_ ( .A(_33_ ), .Z(\SEG0[1] ) );
BUF_X1 _63_ ( .A(_33_ ), .Z(\SEG0[2] ) );
BUF_X1 _64_ ( .A(_33_ ), .Z(\SEG0[3] ) );
BUF_X1 _65_ ( .A(_33_ ), .Z(\SEG0[4] ) );
BUF_X1 _66_ ( .A(_33_ ), .Z(\SEG0[5] ) );
BUF_X1 _67_ ( .A(_33_ ), .Z(\SEG0[6] ) );
BUF_X1 _68_ ( .A(_33_ ), .Z(\SEG0[7] ) );
BUF_X1 _69_ ( .A(\SW[6] ), .Z(_16_ ) );
BUF_X1 _70_ ( .A(\SW[7] ), .Z(_17_ ) );
BUF_X1 _71_ ( .A(\SW[5] ), .Z(_15_ ) );
BUF_X1 _72_ ( .A(\SW[4] ), .Z(_14_ ) );
BUF_X1 _73_ ( .A(\SW[3] ), .Z(_13_ ) );
BUF_X1 _74_ ( .A(\SW[2] ), .Z(_12_ ) );
BUF_X1 _75_ ( .A(\SW[1] ), .Z(_11_ ) );
BUF_X1 _76_ ( .A(_00_ ), .Z(LD4 ) );
BUF_X1 _77_ ( .A(_03_ ), .Z(\LD[2] ) );
BUF_X1 _78_ ( .A(_02_ ), .Z(\LD[1] ) );
BUF_X1 _79_ ( .A(_01_ ), .Z(\LD[0] ) );
BUF_X1 _80_ ( .A(_08_ ), .Z(\SEG[4] ) );
BUF_X1 _81_ ( .A(_06_ ), .Z(\SEG[2] ) );
BUF_X1 _82_ ( .A(_10_ ), .Z(\SEG[6] ) );
BUF_X1 _83_ ( .A(_09_ ), .Z(\SEG[5] ) );
BUF_X1 _84_ ( .A(_07_ ), .Z(\SEG[3] ) );
BUF_X1 _85_ ( .A(_05_ ), .Z(\SEG[1] ) );
BUF_X1 _86_ ( .A(_04_ ), .Z(\SEG[0] ) );

endmodule
