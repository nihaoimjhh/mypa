//Generate the verilog at 2024-08-20T00:45:00
module top (
clk,
reset,
hex_high,
hex_low,
out
);

input clk ;
input reset ;
output [6:0] hex_high ;
output [6:0] hex_low ;
output [7:0] out ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire clk ;
wire reset ;
wire x8 ;
wire [6:0] hex_high ;
wire [6:0] hex_low ;
wire [7:0] out ;


AND2_X1 _092_ ( .A1(_076_ ), .A2(_075_ ), .ZN(_024_ ) );
INV_X1 _093_ ( .A(_077_ ), .ZN(_025_ ) );
NOR2_X1 _094_ ( .A1(_024_ ), .A2(_025_ ), .ZN(_026_ ) );
INV_X1 _095_ ( .A(_026_ ), .ZN(_027_ ) );
INV_X1 _096_ ( .A(_078_ ), .ZN(_028_ ) );
OAI211_X2 _097_ ( .A(_027_ ), .B(_028_ ), .C1(_004_ ), .C2(_077_ ), .ZN(_029_ ) );
OR4_X4 _098_ ( .A1(_076_ ), .A2(_028_ ), .A3(_075_ ), .A4(_005_ ), .ZN(_030_ ) );
NAND2_X1 _099_ ( .A1(_029_ ), .A2(_030_ ), .ZN(_017_ ) );
INV_X1 _100_ ( .A(_076_ ), .ZN(_031_ ) );
NAND4_X1 _101_ ( .A1(_031_ ), .A2(_075_ ), .A3(_077_ ), .A4(_078_ ), .ZN(_032_ ) );
OAI21_X1 _102_ ( .A(_028_ ), .B1(_076_ ), .B2(_075_ ), .ZN(_033_ ) );
OAI21_X1 _103_ ( .A(_032_ ), .B1(_026_ ), .B2(_033_ ), .ZN(_018_ ) );
NAND4_X1 _104_ ( .A1(_031_ ), .A2(_075_ ), .A3(_005_ ), .A4(_078_ ), .ZN(_034_ ) );
AOI21_X1 _105_ ( .A(_075_ ), .B1(_031_ ), .B2(_077_ ), .ZN(_035_ ) );
OAI21_X1 _106_ ( .A(_034_ ), .B1(_035_ ), .B2(_078_ ), .ZN(_019_ ) );
INV_X1 _107_ ( .A(_075_ ), .ZN(_036_ ) );
NOR2_X1 _108_ ( .A1(_036_ ), .A2(_076_ ), .ZN(_037_ ) );
AOI21_X1 _109_ ( .A(_078_ ), .B1(_037_ ), .B2(_025_ ), .ZN(_038_ ) );
NAND3_X1 _110_ ( .A1(_031_ ), .A2(_036_ ), .A3(_077_ ), .ZN(_039_ ) );
NOR3_X1 _111_ ( .A1(_031_ ), .A2(_075_ ), .A3(_077_ ), .ZN(_040_ ) );
INV_X1 _112_ ( .A(_040_ ), .ZN(_041_ ) );
AOI22_X1 _113_ ( .A1(_038_ ), .A2(_039_ ), .B1(_041_ ), .B2(_078_ ), .ZN(_042_ ) );
AND2_X1 _114_ ( .A1(_024_ ), .A2(_077_ ), .ZN(_043_ ) );
OR2_X1 _115_ ( .A1(_042_ ), .A2(_043_ ), .ZN(_020_ ) );
OAI211_X2 _116_ ( .A(_077_ ), .B(_078_ ), .C1(_036_ ), .C2(_076_ ), .ZN(_044_ ) );
OAI21_X1 _117_ ( .A(_044_ ), .B1(_041_ ), .B2(_078_ ), .ZN(_021_ ) );
MUX2_X1 _118_ ( .A(_025_ ), .B(_031_ ), .S(_075_ ), .Z(_045_ ) );
OAI22_X1 _119_ ( .A1(_027_ ), .A2(_033_ ), .B1(_045_ ), .B2(_028_ ), .ZN(_022_ ) );
AND3_X1 _120_ ( .A1(_031_ ), .A2(_075_ ), .A3(_077_ ), .ZN(_046_ ) );
AOI21_X1 _121_ ( .A(_046_ ), .B1(_025_ ), .B2(_024_ ), .ZN(_047_ ) );
AOI22_X1 _122_ ( .A1(_047_ ), .A2(_078_ ), .B1(_038_ ), .B2(_039_ ), .ZN(_023_ ) );
INV_X1 _123_ ( .A(_082_ ), .ZN(_048_ ) );
OR4_X4 _124_ ( .A1(_080_ ), .A2(_048_ ), .A3(_079_ ), .A4(_006_ ), .ZN(_049_ ) );
AND2_X1 _125_ ( .A1(_080_ ), .A2(_079_ ), .ZN(_050_ ) );
AND2_X1 _126_ ( .A1(_050_ ), .A2(_081_ ), .ZN(_051_ ) );
INV_X1 _127_ ( .A(_081_ ), .ZN(_052_ ) );
AOI21_X1 _128_ ( .A(_051_ ), .B1(_007_ ), .B2(_052_ ), .ZN(_053_ ) );
OAI21_X1 _129_ ( .A(_049_ ), .B1(_053_ ), .B2(_082_ ), .ZN(_010_ ) );
INV_X1 _130_ ( .A(_080_ ), .ZN(_054_ ) );
NAND4_X1 _131_ ( .A1(_054_ ), .A2(_079_ ), .A3(_081_ ), .A4(_082_ ), .ZN(_055_ ) );
NOR2_X1 _132_ ( .A1(_050_ ), .A2(_052_ ), .ZN(_056_ ) );
OAI21_X1 _133_ ( .A(_048_ ), .B1(_080_ ), .B2(_079_ ), .ZN(_057_ ) );
OAI21_X1 _134_ ( .A(_055_ ), .B1(_056_ ), .B2(_057_ ), .ZN(_011_ ) );
NAND4_X1 _135_ ( .A1(_054_ ), .A2(_079_ ), .A3(_006_ ), .A4(_082_ ), .ZN(_058_ ) );
AOI21_X1 _136_ ( .A(_079_ ), .B1(_054_ ), .B2(_081_ ), .ZN(_059_ ) );
OAI21_X1 _137_ ( .A(_058_ ), .B1(_059_ ), .B2(_082_ ), .ZN(_012_ ) );
INV_X1 _138_ ( .A(_079_ ), .ZN(_060_ ) );
NOR2_X1 _139_ ( .A1(_060_ ), .A2(_080_ ), .ZN(_061_ ) );
AOI21_X1 _140_ ( .A(_082_ ), .B1(_061_ ), .B2(_052_ ), .ZN(_062_ ) );
NAND3_X1 _141_ ( .A1(_054_ ), .A2(_060_ ), .A3(_081_ ), .ZN(_063_ ) );
NOR3_X1 _142_ ( .A1(_054_ ), .A2(_079_ ), .A3(_081_ ), .ZN(_064_ ) );
INV_X1 _143_ ( .A(_064_ ), .ZN(_065_ ) );
AOI22_X1 _144_ ( .A1(_062_ ), .A2(_063_ ), .B1(_065_ ), .B2(_082_ ), .ZN(_066_ ) );
OR2_X1 _145_ ( .A1(_066_ ), .A2(_051_ ), .ZN(_013_ ) );
OAI211_X2 _146_ ( .A(_081_ ), .B(_082_ ), .C1(_060_ ), .C2(_080_ ), .ZN(_067_ ) );
OAI21_X1 _147_ ( .A(_067_ ), .B1(_065_ ), .B2(_082_ ), .ZN(_014_ ) );
OR3_X2 _148_ ( .A1(_057_ ), .A2(_050_ ), .A3(_052_ ), .ZN(_068_ ) );
MUX2_X1 _149_ ( .A(_052_ ), .B(_054_ ), .S(_079_ ), .Z(_069_ ) );
OAI21_X1 _150_ ( .A(_068_ ), .B1(_048_ ), .B2(_069_ ), .ZN(_015_ ) );
AND3_X1 _151_ ( .A1(_054_ ), .A2(_079_ ), .A3(_081_ ), .ZN(_070_ ) );
AOI21_X1 _152_ ( .A(_070_ ), .B1(_052_ ), .B2(_050_ ), .ZN(_071_ ) );
AOI22_X1 _153_ ( .A1(_071_ ), .A2(_082_ ), .B1(_062_ ), .B2(_063_ ), .ZN(_016_ ) );
INV_X1 _154_ ( .A(_083_ ), .ZN(_008_ ) );
XNOR2_X2 _155_ ( .A(_078_ ), .B(_079_ ), .ZN(_072_ ) );
XNOR2_X2 _156_ ( .A(_075_ ), .B(_005_ ), .ZN(_073_ ) );
XNOR2_X1 _157_ ( .A(_072_ ), .B(_073_ ), .ZN(_074_ ) );
MUX2_X2 _158_ ( .A(_084_ ), .B(_074_ ), .S(_008_ ), .Z(_009_ ) );
DFF_X1 _159_ ( .D(_091_ ), .CK(clk ), .Q(x8 ), .QN(_089_ ) );
DFFS_X1 _160_ ( .D(\out [1] ), .SN(_090_ ), .CK(clk ), .Q(\out [0] ), .QN(_088_ ) );
DFFR_X1 _161_ ( .D(\out [2] ), .RN(_090_ ), .CK(clk ), .Q(\out [1] ), .QN(_000_ ) );
DFFR_X1 _162_ ( .D(\out [3] ), .RN(_090_ ), .CK(clk ), .Q(\out [2] ), .QN(_001_ ) );
DFFR_X1 _163_ ( .D(\out [4] ), .RN(_090_ ), .CK(clk ), .Q(\out [3] ), .QN(_087_ ) );
DFFR_X1 _164_ ( .D(\out [5] ), .RN(_090_ ), .CK(clk ), .Q(\out [4] ), .QN(_086_ ) );
DFFR_X1 _165_ ( .D(\out [6] ), .RN(_090_ ), .CK(clk ), .Q(\out [5] ), .QN(_003_ ) );
DFFR_X1 _166_ ( .D(\out [7] ), .RN(_090_ ), .CK(clk ), .Q(\out [6] ), .QN(_002_ ) );
DFFR_X1 _167_ ( .D(x8 ), .RN(_090_ ), .CK(clk ), .Q(\out [7] ), .QN(_085_ ) );
BUF_X1 _168_ ( .A(\out [1] ), .Z(_076_ ) );
BUF_X1 _169_ ( .A(\out [0] ), .Z(_075_ ) );
BUF_X1 _170_ ( .A(_000_ ), .Z(_004_ ) );
BUF_X1 _171_ ( .A(\out [2] ), .Z(_077_ ) );
BUF_X1 _172_ ( .A(_001_ ), .Z(_005_ ) );
BUF_X1 _173_ ( .A(\out [3] ), .Z(_078_ ) );
BUF_X1 _174_ ( .A(_017_ ), .Z(\hex_low [0] ) );
BUF_X1 _175_ ( .A(_018_ ), .Z(\hex_low [1] ) );
BUF_X1 _176_ ( .A(_019_ ), .Z(\hex_low [2] ) );
BUF_X1 _177_ ( .A(_020_ ), .Z(\hex_low [3] ) );
BUF_X1 _178_ ( .A(_021_ ), .Z(\hex_low [4] ) );
BUF_X1 _179_ ( .A(_022_ ), .Z(\hex_low [5] ) );
BUF_X1 _180_ ( .A(_023_ ), .Z(\hex_low [6] ) );
BUF_X1 _181_ ( .A(\out [5] ), .Z(_080_ ) );
BUF_X1 _182_ ( .A(\out [4] ), .Z(_079_ ) );
BUF_X1 _183_ ( .A(_003_ ), .Z(_007_ ) );
BUF_X1 _184_ ( .A(\out [6] ), .Z(_081_ ) );
BUF_X1 _185_ ( .A(_002_ ), .Z(_006_ ) );
BUF_X1 _186_ ( .A(\out [7] ), .Z(_082_ ) );
BUF_X1 _187_ ( .A(_010_ ), .Z(\hex_high [0] ) );
BUF_X1 _188_ ( .A(_011_ ), .Z(\hex_high [1] ) );
BUF_X1 _189_ ( .A(_012_ ), .Z(\hex_high [2] ) );
BUF_X1 _190_ ( .A(_013_ ), .Z(\hex_high [3] ) );
BUF_X1 _191_ ( .A(_014_ ), .Z(\hex_high [4] ) );
BUF_X1 _192_ ( .A(_015_ ), .Z(\hex_high [5] ) );
BUF_X1 _193_ ( .A(_016_ ), .Z(\hex_high [6] ) );
BUF_X1 _194_ ( .A(reset ), .Z(_083_ ) );
BUF_X1 _195_ ( .A(_008_ ), .Z(_090_ ) );
BUF_X1 _196_ ( .A(x8 ), .Z(_084_ ) );
BUF_X1 _197_ ( .A(_009_ ), .Z(_091_ ) );

endmodule
